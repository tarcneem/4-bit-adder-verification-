module adder(
    input [3:0] A,B,
    output [4:0] Y
        );
      
    assign Y = A + B;  
      
    endmodule